  module multiplier_8bit
  ( input [7:0] A,B,
   output [7:0] P );
  assign P = A*B;
endmodule
  